----------------------------------------------------------------------------------
-- FPGA Design Using VHDL
-- Final Project
--
-- Authors: Eric Beales &  James Frank
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

package final_project_lib is

type byte_array is array (integer range <>) of unsigned(7 downto 0);

end final_project_lib;

package body final_project_lib is
 
end final_project_lib;
